module fn_menor (
    output Y,
    input  a,
    input  b
);
    assign Y = a & b;
endmodule
