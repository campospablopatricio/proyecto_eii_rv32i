//Función *MENOR QUE* de 32 bit para valores en binario natural y con signo complemento a dos. Incluye 
//una entrada de selección, $0$ con signo y $1$ sin signo, dos entradas, $A$ y $B$, de 32 bit y una 
//salida de un bit. 
//La salida es $1$ si la entrada $A$ es menor que la entrada $B$ y $0$ caso contrario. 
//La comparación se realiza considerando valores en binario natural o en complemento a dos según indique 
//la entrada de selección.
  
module fn_menor (
    input  [31 : 0] a,
    input  [31 : 0] b,
    input           sin_signo,
    output          Y
);
 
  assign Y = sin_signo ? (a < b) : ($signed(a) < $signed(b));
  
endmodule

//otra forma de hacerlo, sin usar signed (propio de verilog), 
//es con el bit mas significativo de a y b osea a[31] y b[31] 
//con signo para 0 y 1 caso contrario. 1 si a<b y 0 si b<a
