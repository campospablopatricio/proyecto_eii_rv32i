module and1 (
    output Y,
    input  a,
    input  b
);
    assign Y = a & b;
endmodule
